
`define MAX_DUTY 1000000
`define MIN_DUTY 1
`define DUTY_STEP 1000
`define REG_LEN 20
// Two debounced buttons are used to control the duty cycle (step size: 10%)
module PWM_Generator_Verilog
 (
    clk, // 100MHz clock input 
    duty_val,
    val_en,
    increase_duty, // input to increase 10% duty cycle 
    decrease_duty, // input to decrease 10% duty cycle 
    PWM_OUT // 10MHz PWM output signal 
);

initial begin
    $dumpfile("pwm.vcd");
    $dumpvars(0, PWM_Generator_Verilog);
end
 input clk;
 input [`REG_LEN:0]duty_val;
 input val_en;
 input increase_duty;
 input decrease_duty;
 output PWM_OUT;
 wire slow_clk_enable; // slow clock enable signal for debouncing FFs
 reg[27:0] counter_debounce=0;// counter for creating slow clock enable signals 
 reg [31:0]counter=0;

 wire tmp1,tmp2,duty_inc;// temporary flip-flop signals for debouncing the increasing button
 wire tmp3,tmp4,duty_dec;// temporary flip-flop signals for debouncing the decreasing button
 reg[`REG_LEN:0] counter_PWM=0;// counter for creating 10Mhz PWM signal
 reg[`REG_LEN:0] DUTY_CYCLE=`MAX_DUTY / 2; // initial duty cycle is 50%
  // Debouncing 2 buttons for inc/dec duty cycle 
  // Firstly generate slow clock enable for debouncing flip-flop (4Hz)

 always @(posedge clk) begin
    counter <= counter + 1;
    if (counter[4:0] === 0) 
        $display("%d", counter);
    if (counter > 10000000)
        $finish;
    counter_debounce <= counter_debounce + 1;
    //if(counter_debounce>=25000000) then  
    // for running on FPGA -- comment when running simulation
    if(counter_debounce>=1) 
    // for running simulation -- comment when running on FPGA
        counter_debounce <= 0;
    end
 // assign slow_clk_enable = counter_debounce == 25000000 ?1:0;
 // for running on FPGA -- comment when running simulation 
 assign slow_clk_enable = counter_debounce == 1 ?1:0;
 // for running simulation -- comment when running on FPGA
 // debouncing FFs for increasing button
 DFF_PWM PWM_DFF1(clk,slow_clk_enable,increase_duty,tmp1);
 DFF_PWM PWM_DFF2(clk,slow_clk_enable,tmp1, tmp2); 
 assign duty_inc =  tmp1 & (~ tmp2) & slow_clk_enable;
 // debouncing FFs for decreasing button
 DFF_PWM PWM_DFF3(clk,slow_clk_enable,decrease_duty, tmp3);
 DFF_PWM PWM_DFF4(clk,slow_clk_enable,tmp3, tmp4); 
 assign duty_dec =  tmp3 & (~ tmp4) & slow_clk_enable;
 // vary the duty cycle using the debounced buttons above
 always @(posedge clk)
    begin
    if (val_en)
        DUTY_CYCLE <= duty_val;
    else if(duty_inc==1 && DUTY_CYCLE <= `MAX_DUTY) 
        DUTY_CYCLE <= DUTY_CYCLE + `DUTY_STEP;// increase duty cycle by 1%
    else if(duty_dec == 1 && DUTY_CYCLE >= `MIN_DUTY + `DUTY_STEP) 
        DUTY_CYCLE <= DUTY_CYCLE - `DUTY_STEP;//decrease duty cycle by 1%
    end 
// Create 10MHz PWM signal with variable duty cycle controlled by 2 buttons 
 always @(posedge clk)
    begin
    counter_PWM <= counter_PWM + 1;
    if(counter_PWM >= `MAX_DUTY) 
        counter_PWM <= 0;
    end
 assign PWM_OUT = counter_PWM < DUTY_CYCLE ? 1:0;
endmodule
// Debouncing DFFs for push buttons on FPGA
module DFF_PWM(clk,en,D,Q);
    input clk,en,D;
    output reg Q;
    always @(posedge clk)
        begin 
            if(en==1) // slow clock enable signal 
            Q <= D;
        end 
endmodule 